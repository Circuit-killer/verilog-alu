module InstructionMemory(
  input [31:0] Address,
  input Clk,
  output reg [31:0] ReadData
);
  parameter NUM_CELLS = 32 - 1;
  reg [31:0] tab[NUM_CELLS:0];

  integer i;
  initial begin
    // Zero all the cells.
    for (i = 0; i <= NUM_CELLS; i = i + 1)
      tab[i] <= 0;

    // addi $1, $0, 1
    tab[0] <= 'b 001000_00000_00001_0000_0000_0000_0001;
    // addi $20, $0, 0xDEAD
    tab[1] <= 'b 001000_00000_10100_1101_1110_1010_1101;
    // sw $20, 0($1)
    tab[2] <= 'b 101011_00001_10100_0000_0000_0000_0000;
    // sw $20, 1($1)
    tab[3] <= 'b 101011_00001_10100_0000_0000_0000_0001;
    // sw $20, 3($0)
    tab[4] <= 'b 101011_00000_10100_0000_0000_0000_0011;

    // add $1, $1, $1
    tab[5] <= 'b 000000_00001_00001_00001_00000_100000;
    // add $1, $1, $1
    tab[6] <= 'b 000000_00001_00001_00001_00000_100000;
    // add $1, $1, $1
    tab[7] <= 'b 000000_00001_00001_00001_00000_100000;

    // lw $4, 1($0)
    tab[8] <= 'b 100011_00000_00100_0000_0000_0000_0011;
    // and $4, $1, $4
    tab[9] <= 'b 000000_00001_00100_00100_00000_100100;

    // j 16
    tab[10] <= 'b 000010_0000_0000_0000_0000_0000_010000;
    // addi $1, $0, 1 (shouldn't be executed)
    tab[11] <= 'b 001000_00000_00001_0000_0000_0000_0001;

    // addi $2, $2, 2
    tab[16] <= 'b 001000_00010_00010_0000_0000_0000_0010;
    // bne $2, $4, -3 (16)
    tab[17] <= 'b 000101_00010_00100_1111_1111_1111_1101;
    // sw $2, 8($0)
    tab[18] <= 'b 101011_00000_00010_0000_0000_0000_1000;
  end

  always @(posedge Clk) begin
    ReadData <= tab[Address];
  end
endmodule
